//======================================================================
//
// chacha_qr.v
// -----------
// Verilog 2001 implementation of the stream cipher ChaCha.
// This is the combinational QR logic as a separade module to allow
// us to build versions of the cipher with 1, 2, 4 and even 8
// parallel qr functions.
//
//
// Copyright (c) 2013 Secworks Sweden AB
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or
// without modification, are permitted provided that the following
// conditions are met:
//
// 1. Redistributions of source code must retain the above copyright
//    notice, this list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright
//    notice, this list of conditions and the following disclaimer in
//    the documentation and/or other materials provided with the
//    distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
// FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
// COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,
// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
// BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
// ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//======================================================================

module chacha_qr(
                 input wire [31 : 0]  a,    //Defining Inputs
                 input wire [31 : 0]  b,
                 input wire [31 : 0]  c,
                 input wire [31 : 0]  d,

                 output wire [31 : 0] a_prim,   //Defining Outputs
                 output wire [31 : 0] b_prim,
                 output wire [31 : 0] c_prim,
                 output wire [31 : 0] d_prim
                );

  //----------------------------------------------------------------
  // Declaring wires for output
  //----------------------------------------------------------------
  reg [31 : 0] internal_a_prim;
  reg [31 : 0] internal_b_prim;
  reg [31 : 0] internal_c_prim;
  reg [31 : 0] internal_d_prim;


  //----------------------------------------------------------------
  // Concurrent connectivity of output ports.
  //----------------------------------------------------------------
  assign a_prim = internal_a_prim;
  assign b_prim = internal_b_prim;
  assign c_prim = internal_c_prim;
  assign d_prim = internal_d_prim;


  //----------------------------------------------------------------
  // qr
  // The actual quarterround function.
  //----------------------------------------------------------------
  always @*
    begin : qr
      reg [31 : 0] a0;                  // Declaring registers for intermediate results
      reg [31 : 0] a1;

      reg [31 : 0] b0;
      reg [31 : 0] b1;                  // Declaring registers for intermediate results
      reg [31 : 0] b2;
      reg [31 : 0] b3;

      reg [31 : 0] c0;
      reg [31 : 0] c1;                  // Declaring registers for intermediate results

      reg [31 : 0] d0;
      reg [31 : 0] d1;                  // Declaring registers for intermediate results
      reg [31 : 0] d2;
      reg [31 : 0] d3;

      a0 = a + b;                       // First Step of Quarterround : 32 bit addition
      d0 = d ^ a0;                      // Second Step of Quarterround : 32 bit XOR Operation
      d1 = {d0[15 : 0], d0[31 : 16]};   // Third Step of Quarterround : Left shifting the bits by 16 bit
      
      c0 = c + d1;                       // First Step of Quarterround : 32 bit addition
      b0 = b ^ c0;                       // Second Step of Quarterround : 32 bit XOR Operation
      b1 = {b0[19 : 0], b0[31 : 20]};    // Third Step of Quarterround : Left shifting the bits by 12 bit
      
      a1 = a0 + b1;                      // First Step of Quarterround : 32 bit addition
      d2 = d1 ^ a1;                      // Second Step of Quarterround : 32 bit XOR Operation
      d3 = {d2[23 : 0], d2[31 : 24]};;   // Third Step of Quarterround : Left shifting the bits by 8 bit
     
      c1 = c0 + d3;                      // First Step of Quarterround : 32 bit addition
      b2 = b1 ^ c1;                      // Second Step of Quarterround : 32 bit XOR Operation
      b3 = {b2[24 : 0], b2[31 : 25]};    // Third Step of Quarterround : Left shifting the bits by 7 bit

      internal_a_prim = a1;              // Sequentially connecting output port wires to the intermediate registers 
      internal_b_prim = b3;
      internal_c_prim = c1;
      internal_d_prim = d3;
    end // qr
endmodule // chacha_qr

//======================================================================
// EOF chacha_qr.v
//======================================================================
